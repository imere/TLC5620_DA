module Convert (
	input clk,
	input [3:0] i,      // 2^4 === 16 > 10
	output reg [7:0] o
);

	always @ (posedge clk)
		begin

			case (i)
				// h~a : 0
				8'd0: o <= 8'b11000000;
				8'd1: o <= 8'b11111001;
				8'd2: o <= 8'b10100100;
				8'd3: o <= 8'b10110000;
				8'd4: o <= 8'b10011001;
				8'd5: o <= 8'b10010010;
				8'd6: o <= 8'b10000010;
				8'd7: o <= 8'b11111000;
				8'd8: o <= 8'b10000000;
				8'd9: o <= 8'b10010000;
				8'd10: o <= 8'b10001000;
				8'd11: o <= 8'b10000011;
				8'd12: o <= 8'b11000110;
				8'd13: o <= 8'b10100001;
				8'd14: o <= 8'b10000110;
				8'd15: o <= 8'b10001110;
				default: o <= 8'b10111111;
			endcase

		end

endmodule
